module moduleName (
    input addr[7:0],
    output reg [7:0]
);

always @(posedge clk ) begin
    
end
    
endmodule